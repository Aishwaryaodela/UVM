
	/////////////////////////////////////////////////////////////////////////////////
	//     IN THIS SLAVE SEQUNCER CLASS WE HAVE TO CREATE A CONSTRUCTOR FOR IT     //
	/////////////////////////////////////////////////////////////////////////////////

class apb_slave_sequencer extends uvm_sequencer#(sequence_item);

	`uvm_component_utils(apb_slave_sequencer)     				//------ FACTORY REGISTRATION

	
	//////////////////////////////////////////////////////////////////////////////
	//   NEW CONSTRUCTOR FOR FOR CREATING MEMORY AND POINTING TO THE PARENT     //
	//////////////////////////////////////////////////////////////////////////////

	function new(string name = "apb_slave_sequencer",uvm_component parent);
		super.new(name,parent);
	endfunction

endclass
