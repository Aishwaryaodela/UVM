
	//////////////////////////////////////////////////////////////////////////////////
	//     IN THIS MASTER SEQUNCER CLASS WE HAVE TO CREATE A CONSTRUCTOR FOR IT     //
	//////////////////////////////////////////////////////////////////////////////////

class master_sequencer extends uvm_sequencer#(sequence_item);

	`uvm_component_utils(master_sequencer)     					//------ FACTORY REGISTRATION

	
	//////////////////////////////////////////////////////////////////////////////
	//   NEW CONSTRUCTOR FOR FOR CREATING MEMORY AND POINTING TO THE PARENT     //
	//////////////////////////////////////////////////////////////////////////////

	function new(string name = "master_sequencer",uvm_component parent);
		super.new(name,parent);
	endfunction

endclass
