
	//////////////////////////////////////////////////////////////////////////////////
	//     IN THIS RX MAC SEQUNCER CLASS WE HAVE TO CREATE A CONSTRUCTOR FOR IT     //
	//////////////////////////////////////////////////////////////////////////////////

class rx_mac_sequencer extends uvm_sequencer#(sequence_item);

	`uvm_component_utils(rx_mac_sequencer)     						//------ FACTORY REGISTRATION

	
	//////////////////////////////////////////////////////////////////////////////
	//   NEW CONSTRUCTOR FOR FOR CREATING MEMORY AND POINTING TO THE PARENT     //
	//////////////////////////////////////////////////////////////////////////////

	function new(string name = "rx_mac_sequencer",uvm_component parent);
		super.new(name,parent);
	endfunction

endclass
